interface axi_if;

  // clock and reset
  logic clk;
  logic reset_n;

endinterface