class axi_txn;

  logic [31:0] addr;
  logic [31:0] data;
  logic        write;

endclass
